library IEEE;
use IEEE.std_logic_1164.all;

package common is
--    impure function init_mem(input_file : in string) return 
end;

--package body common is
--end common;
